module and_gate(A, B, C);
    input A, B;
    output C;
 
    and(C, A, B);
endmodule